-- Praktikum EL3111 Arsitektur Sistem Komputer
-- Modul : 5
-- Percobaan : 1
-- Tanggal : 1 Desember 2014
-- Kelompok : III
-- Rombongan : A
-- Nama (NIM) 1 : Damon Prasetyo Arso (13212001)
-- Nama (NIM) 2 : Muhammad Mustadi (13210056)
-- Nama File : data_memory.vhd
-- Deskripsi : Program Data Memory


LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY altera_mf;
USE altera_mf.all;
ENTITY data_memory IS
PORT (
ADDR : IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- alamat
WR_EN : IN STD_LOGIC; --Indikator Penulisan
RD_EN : IN STD_LOGIC; --Indikator Pembacaan
clock : IN STD_LOGIC := '1'; -- clock
RD_Data : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
WR_DATA : IN STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE structural of data_memory IS
SIGNAL sub_wire0 : STD_LOGIC_VECTOR (7 DOWNTO 0);
COMPONENT altsyncram
-- komponen memori
GENERIC
(
init_file : STRING; -- name of the .mif file
operation_mode : STRING; -- the operation mode
widthad_a : NATURAL; -- width of address_a[]
width_a : NATURAL -- width of data_a[]
);
PORT
(
wren_a : IN STD_LOGIC; -- Write Enable Activation
clock0 : IN STD_LOGIC ; -- Clock
address_a : IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- Address Input
q_a : OUT STD_LOGIC_VECTOR (7 DOWNTO 0); -- Data Output
data_a : IN STD_LOGIC_VECTOR (7 DOWNTO 0) -- Data Input
);
END COMPONENT;

BEGIN
altsyncram_component : altsyncram
GENERIC MAP
(
init_file => "dmemory.mif",
operation_mode => "SINGLE_PORT",
widthad_a => 8,
width_a => 8
)
PORT MAP
(
wren_a => WR_EN AND NOT RD_EN, -- isi yang sesuai
clock0 => clock,
address_a => ADDR,
q_a => RD_DATA, -- isi yang sesuai
data_a => WR_Data
);

END structural;
