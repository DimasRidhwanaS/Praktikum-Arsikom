-- Praktikum EL3111 Arsitektur Sistem Komputer
-- Modul : 3
-- Percobaan : 4
-- Tanggal : 27 Oktober 2023
-- Kelompok : 2
-- Rombongan : D
-- Nama (NIM) 1 : Dimas Ridhwana Shalsareza (13221076)
-- Nama (NIM) 2 : M. Zhafran Arrafi Anwar (13221079)


LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
LIBRARY altera_mf;
USE altera_mf.all;

ENTITY reg_file IS
	PORT (
		clock : IN STD_LOGIC; -- clock
		WR_EN : IN STD_LOGIC; -- write enable
		ADDR_1 : IN STD_LOGIC_VECTOR (4 DOWNTO 0); -- Input 1
		ADDR_2 : IN STD_LOGIC_VECTOR (4 DOWNTO 0); -- Input 2
		ADDR_3 : IN STD_LOGIC_VECTOR (4 DOWNTO 0); -- Input 3
		WR_Data_3 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);-- write data
		RD_Data_1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);-- read data 1
		RD_Data_2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) -- read data 2
		);
END ENTITY;

ARCHITECTURE behavior OF reg_file IS
TYPE ramtype IS ARRAY (31 DOWNTO 0) OF std_logic_vector (31 DOWNTO 0);
SIGNAL mem: ramtype;
	BEGIN
		PROCESS (clock, WR_EN, ADDR_1, ADDR_2, ADDR_3)
		BEGIN
			IF ((clock'EVENT) and (clock = '0') and WR_EN = '0') THEN
				RD_Data_1 <= mem(conv_integer((ADDR_1)));
				RD_Data_2 <= mem(conv_integer((ADDR_2)));
			ELSIF ((clock'EVENT) and (clock = '1') and WR_EN = '1') THEN
				mem(conv_integer((ADDR_3))) <= WR_Data_3;
			END IF;
		END PROCESS;
END behavior;