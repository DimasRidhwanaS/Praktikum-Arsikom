LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY bus_merger IS
PORT (
    DATA_IN1 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    DATA_IN2 : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
    DATA_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
);
END bus_merger;

ARCHITECTURE arch_bus_merger OF bus_merger IS
BEGIN
    DATA_OUT <= DATA_IN2 & DATA_IN1;
END arch_bus_merger;