-- Praktikum EL3111 Arsitektur Sistem Komputer
-- Modul : 5
-- Percobaan : 1
-- Tanggal : 1 Desember 2014
-- Kelompok : III
-- Rombongan : A
-- Nama (NIM) 1 : Damon Prasetyo Arso (13212001)
-- Nama (NIM) 2 : Muhammad Mustadi (13210056)
-- Nama File : comparator.vhd
-- Deskripsi : Program Comparator

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY comparator IS
  PORT (
    D_1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    D_2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    EQ : OUT STD_LOGIC -- Hasil Perbandingan EQ
  );
END comparator;

ARCHITECTURE comp OF comparator IS
  BEGIN
  PROCESS (D_1,D_2)
		BEGIN
			IF (D_1 = D_2) THEN
				EQ <= '1';
			ELSE 
				EQ <= '0';
			END IF;
		END PROCESS;
  END comp;